`timescale 1ns / 1ps
module alu_tb;

	// Inputs
	reg [31:0] A;
	reg [31:0] B;
	reg [3:0] Op;

	// Outputs
	wire [31:0] Out;
	wire Zero;

	// Instantiate the Unit Under Test (UUT)
	alu uut (
		.Out(Out), 
		.Zero(Zero), 
		.A(A), 
		.B(B), 
		.Op(Op)
	);

	initial begin
		// Initialize Inputs
		A = 32'b00000000000000000000000000000001;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b0000;
		#5;
		
		A = 32'b00000000000000000000000000000010;
		B = 32'b00000000000000000000000000000001;
		Op = 4'b0001;
		#5;
		
		A = 32'b00000000000000000000000000000011;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b0010;
		#5;

		A = 32'b00000000000000000000000000000001;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b0011;
		#5;

		A = 32'b00000000000000000000000000000001;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b0100;
		#5;
		
		A = 32'b11111111111111111111111111111111;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b1000;
		#5;
		
		A = 32'b00111111111111111111111111111111;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b1000;
		#5;
		
		A = 32'b00111111111111111111111111111111;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b1010;
		#5;
		
		A = 32'b11111111111111111111111111111111;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b1010;
		#5;
		
		A = 32'b11111111111111111111111111111110;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b1000;
		#5;


 		A = 32'b10000011111111111111111111111111;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b1100;
		#5;

 		A = 32'b10000011111111111111111111111111;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b1101;
		#5;
		
 		A = 32'b00000000000000000000000000000001;
		B = 32'b00000000000000000000000000000010;
		Op = 4'b1010;
		#5;


	end
      
endmodule
